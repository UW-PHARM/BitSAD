`timescale 1ns / 1ps
/////////////////////////////////////////////////////////////////////////////////////
// PHARM
// Carly Schulz
//
// determ_mult
//		multiplication unit for the deterministic bitstream 1 = 1 and 0 = -1
/////////////////////////////////////////////////////////////////////////////////////
module determ_mult(a, b, y);

// I/O
input a, b;
output y;

assign y = ~(a ^ b);

endmodule